library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity sync_rom_8_bits is
     port(clk : in std_logic;
     addr_r : in std_logic_vector(7 downto 0);
     data : out std_logic_vector(3 downto 0)
     );
end sync_rom_8_bits;

architecture arch of sync_rom_8_bits is
     constant ADDR_WIDTH : integer:=8;
     constant DATA_WIDTH : integer:=4;
     type rom_type is array (0 to 2**ADDR_WIDTH-1)
         of std_logic_vector(DATA_WIDTH-1 downto 0);
 
-- ROM definition
 constant HEX2LED_LOOK_UP_TABLE: rom_type:=( 
    -- 2^16-by-8
    "00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110100",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110101",
"01110100",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01110110",
"01110101",
"01110100",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01110111",
"01110110",
"01110101",
"01110100",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111000",
"01110111",
"01110110",
"01110101",
"01110100",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111001",
"01111000",
"01110111",
"01110110",
"01110101",
"01110100",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111010",
"01111001",
"01111000",
"01110111",
"01110110",
"01110101",
"01110100",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111011",
"01111010",
"01111001",
"01111000",
"01110111",
"01110110",
"01110101",
"01110100",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"10000011",
"01111101",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111100",
"01111011",
"01111010",
"01111001",
"01111000",
"01110111",
"01110110",
"01110101",
"01110100",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"10000010",
"01111110",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111101",
"01111100",
"01111011",
"01111010",
"01111001",
"01111000",
"01110111",
"01110110",
"01110101",
"01110100",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"10000001",
"01111111",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"01111110",
"01111101",
"01111100",
"01111011",
"01111010",
"01111001",
"01111000",
"01110111",
"01110110",
"01110101",
"01110100",
"01110011",
"01110010",
"01110001",
"01110000",
"01101111",
"01101110",
"01101101",
"01101100",
"01101011",
"01101010",
"01101001",
"01101000",
"01100111",
"01100110",
"01100101",
"01100100",
"01100011",
"01100010",
"01100001",
"01100000",
"01011111",
"01011110",
"01011101",
"01011100",
"01011011",
"01011010",
"01011001",
"01011000",
"01010111",
"01010110",
"01010101",
"01010100",
"01010011",
"01010010",
"01010001",
"01010000",
"01001111",
"01001110",
"01001101",
"01001100",
"01001011",
"01001010",
"01001001",
"01001000",
"01000111",
"01000110",
"01000101",
"01000100",
"01000011",
"01000010",
"01000001",
"01000000",
"00111111",
"00111110",
"00111101",
"00111100",
"00111011",
"00111010",
"00111001",
"00111000",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00101111",
"00101110",
"00101101",
"00101100",
"00101011",
"00101010",
"00101001",
"00101000",
"00100111",
"00100110",
"00100101",
"00100100",
"00100011",
"00100010",
"00100001",
"00100000",
"00011111",
"00011110",
"00011101",
"00011100",
"00011011",
"00011010",
"00011001",
"00011000",
"00010111",
"00010110",
"00010101",
"00010100",
"00010011",
"00010010",
"00010001",
"00010000",
"00001111",
"00001110",
"00001101",
"00001100",
"00001011",
"00001010",
"00001001",
"00001000",
"00000111",
"00000110",
"00000101",
"00000100",
"00000011",
"00000010",
"00000001",
"00000000",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"01111111",
"00000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"01111110",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"01111101",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"01111100",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"01111011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"01111010",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"01110011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"01110010",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"01110001",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"01110000",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"01101111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"01101110",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"01101101",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"01101100",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"01101011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01101010",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"01100011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"01100010",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"01100001",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"01100000",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"01011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"01011110",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"01011101",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"01011100",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"01011011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01011010",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"01010011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"01010010",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"01010001",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"01010000",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"01001111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"01001110",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"01001101",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"01001100",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"01001011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01001010",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"01000011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"01000010",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"01000001",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"01000000",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"00111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"00111110",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"00111101",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"00111100",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"00111011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"00111010",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"00110011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"00110010",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"00110001",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"00110000",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"00101111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"00101110",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"00101101",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"00101100",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"00101011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00101010",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"00100011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"00100010",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"00100001",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"00100000",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"00011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"00011110",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"00011101",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"00011100",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"00011011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00011010",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"00010011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"00010010",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"00010001",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"00010000",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"00001111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"00001110",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"00001101",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"00001100",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110100",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"00001011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110101",
"11110100",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00001010",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110110",
"11110101",
"11110100",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110111",
"11110110",
"11110101",
"11110100",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11111000",
"11110111",
"11110110",
"11110101",
"11110100",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111001",
"11111000",
"11110111",
"11110110",
"11110101",
"11110100",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111010",
"11111001",
"11111000",
"11110111",
"11110110",
"11110101",
"11110100",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111011",
"11111010",
"11111001",
"11111000",
"11110111",
"11110110",
"11110101",
"11110100",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"11111011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111100",
"11111011",
"11111010",
"11111001",
"11111000",
"11110111",
"11110110",
"11110101",
"11110100",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"00000011",
"11111100",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111101",
"11111100",
"11111011",
"11111010",
"11111001",
"11111000",
"11110111",
"11110110",
"11110101",
"11110100",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"00000010",
"11111101",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111110",
"11111101",
"11111100",
"11111011",
"11111010",
"11111001",
"11111000",
"11110111",
"11110110",
"11110101",
"11110100",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"00000001",
"11111110",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111111",
"11111110",
"11111101",
"11111100",
"11111011",
"11111010",
"11111001",
"11111000",
"11110111",
"11110110",
"11110101",
"11110100",
"11110011",
"11110010",
"11110001",
"11110000",
"11101111",
"11101110",
"11101101",
"11101100",
"11101011",
"11101010",
"11101001",
"11101000",
"11100111",
"11100110",
"11100101",
"11100100",
"11100011",
"11100010",
"11100001",
"11100000",
"11011111",
"11011110",
"11011101",
"11011100",
"11011011",
"11011010",
"11011001",
"11011000",
"11010111",
"11010110",
"11010101",
"11010100",
"11010011",
"11010010",
"11010001",
"11010000",
"11001111",
"11001110",
"11001101",
"11001100",
"11001011",
"11001010",
"11001001",
"11001000",
"11000111",
"11000110",
"11000101",
"11000100",
"11000011",
"11000010",
"11000001",
"11000000",
"10111111",
"10111110",
"10111101",
"10111100",
"10111011",
"10111010",
"10111001",
"10111000",
"10110111",
"10110110",
"10110101",
"10110100",
"10110011",
"10110010",
"10110001",
"10110000",
"10101111",
"10101110",
"10101101",
"10101100",
"10101011",
"10101010",
"10101001",
"10101000",
"10100111",
"10100110",
"10100101",
"10100100",
"10100011",
"10100010",
"10100001",
"10100000",
"10011111",
"10011110",
"10011101",
"10011100",
"10011011",
"10011010",
"10011001",
"10011000",
"10010111",
"10010110",
"10010101",
"10010100",
"10010011",
"10010010",
"10010001",
"10010000",
"10001111",
"10001110",
"10001101",
"10001100",
"10001011",
"10001010",
"10001001",
"10001000",
"10000111",
"10000110",
"10000101",
"10000100",
"10000011",
"10000010",
"10000001",
"00000000",
"11111111",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10001010",
"10001011",
"10001100",
"10001101",
"10001110",
"10001111",
"10010000",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001",
"10011010",
"10011011",
"10011100",
"10011101",
"10011110",
"10011111",
"10100000",
"10100001",
"10100010",
"10100011",
"10100100",
"10100101",
"10100110",
"10100111",
"10101000",
"10101001",
"10101010",
"10101011",
"10101100",
"10101101",
"10101110",
"10101111",
"10110000",
"10110001",
"10110010",
"10110011",
"10110100",
"10110101",
"10110110",
"10110111",
"10111000",
"10111001",
"10111010",
"10111011",
"10111100",
"10111101",
"10111110",
"10111111",
"11000000",
"11000001",
"11000010",
"11000011",
"11000100",
"11000101",
"11000110",
"11000111",
"11001000",
"11001001",
"11001010",
"11001011",
"11001100",
"11001101",
"11001110",
"11001111",
"11010000",
"11010001",
"11010010",
"11010011",
"11010100",
"11010101",
"11010110",
"11010111",
"11011000",
"11011001",
"11011010",
"11011011",
"11011100",
"11011101",
"11011110",
"11011111",
"11100000",
"11100001",
"11100010",
"11100011",
"11100100",
"11100101",
"11100110",
"11100111",
"11101000",
"11101001",
"11101010",
"11101011",
"11101100",
"11101101",
"11101110",
"11101111",
"11110000",
"11110001",
"11110010",
"11110011",
"11110100",
"11110101",
"11110110",
"11110111",
"11111000",
"11111001",
"11111010",
"11111011",
"11111100",
"11111101",
"11111110"
     );
 signal rom : rom_type := HEX2LED_LOOK_UP_TABLE ;

begin
 process(clk)
     begin
     if (clk'event and clk = '1') then
     data <= rom(to_integer(unsigned(addr_r)));
     end if;
 end process;
end arch;

